v1 1 0 5
r1 1 2 1
c1 2 0 1e-6

