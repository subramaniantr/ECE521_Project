vdd 1 0 5
mp1 2 3 1 1 pmos 20e-6 1e-6
mn1 2 3 0 0 nmos 10e-6 1e-6
cl1 2 0 1e-12
mp2 4 2 1 1 pmos 20e-6 1e-6
mn2 4 2 0 0 nmos 10e-6 1e-6
cl2 4 0 1e-12
mp3 3 4 1 1 pmos 20e-6 1e-6
mn3 3 4 0 0 nmos 10e-6 1e-6
cl3 3 0 1e-12
