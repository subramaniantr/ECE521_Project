v1 1 0 5
c1 1 2 1e-6
r1 2 0 1
