vdd 1 0 5
c1 2 3 25e-12
c2 3 0 100e-12
lm 1 2 12.665e-6
rl 1 2 10e3
vd 2 4 0
m1 4 0 3 3 nmos 10e-6 1e-6
iss 3 5 0.25e-3
vss 5 0 -5
