v1 1 0 5
r2 1 3 1000
r1 1 2 1
c1 2 0 1e-6
c2 3 0 1e-6

