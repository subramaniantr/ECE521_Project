r1 1 2 1000
r2 2 3 500
r3 3 4 300
r4 4 0 200
u1 1 0 1e-12
